library verilog;
use verilog.vl_types.all;
entity ANDtest is
end ANDtest;
