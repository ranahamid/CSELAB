library verilog;
use verilog.vl_types.all;
entity NANDtest is
end NANDtest;
