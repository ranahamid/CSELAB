library verilog;
use verilog.vl_types.all;
entity NOTtest is
end NOTtest;
