library verilog;
use verilog.vl_types.all;
entity NORtest is
end NORtest;
