library verilog;
use verilog.vl_types.all;
entity XORtest is
end XORtest;
