library verilog;
use verilog.vl_types.all;
entity ORtest is
end ORtest;
